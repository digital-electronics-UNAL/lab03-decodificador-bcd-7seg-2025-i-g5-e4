module Lab3 (
    input clk,
    input [7:0] A,   // Ignorados en esta prueba
    input [7:0] B,
    input Sel,
    output [6:0] SSeg,
    output [3:0] an
);

    wire clk_div;
    wire [1:0] sel_disp;
    reg [3:0] bcd;

    // ✅ Divisor de frecuencia
    DivFrec div_clk (
        .clk(clk),
        .clk_out(clk_div)
    );

    // ✅ Selección de display activo
    SelAn seleccion (
        .clk(clk_div),
        .sel(sel_disp),
        .an(an)
    );

    // ✅ Asignar manualmente los valores para mostrar "1234"
    always @(*) begin
        case (sel_disp)
            2'b00: bcd = 4'd4; // unidades → display derecho (4°)
            2'b01: bcd = 4'd1; // signo → display izquierdo (1°)
            2'b10: bcd = 4'd2; // centenas → 2°
            2'b11: bcd = 4'd3; // decenas → 3°
        endcase
    end

    // ✅ Decodificación a 7 segmentos
    BCDtoSSeg seg (
        .BCD(bcd),
        .SSeg(SSeg)
    );

endmodule
